module pipeid(mwreg,mrn,ern,ewreg,em2reg,mm2reg,dpc4,inst,wrn,wdi,ealu,malu,mmo,wwreg,clk,clrn,bpc,jpc,pcsrc,nostall,wreg,m2reg,wmem,aluc,aluimm,a,b,dimm,rn,shift,jal);
input clk, clrn; 
input [31:0] dpc4;
input [31:0] inst;
input [31:0] wdi; 
input [31:0] ealu; 
input [31:0] malu; 
input [31:0] mmo;
input [4:0] ern; 
input [4:0] mrn; 
input [4:0] wrn; 
input ewreg; 
input em2reg;
input mwreg; 
input mm2reg; 
input wwreg; 
output [31:0] bpc; 
output [31:0] jpc; 
output [31:0] a, b; 
output [31:0] dimm; 
output [4:0] rn; 
output [3:0] aluc; 
output [1:0] pcsrc; 
output nostall;
output wreg; 
output m2reg;
output wmem; 
output aluimm; 
output shift;
output jal; 
wire [5:0] op = inst[31:26]; 
wire [4:0] rs = inst[25:21]; 
wire [4:0] rt = inst[20:16]; 
wire [4:0] rd = inst[15:11]; 
wire [5:0] func = inst[05:00]; 
wire [15:0] imm = inst[15:00]; 
wire [25:0] addr = inst[25:00]; 
wire regrt;
wire sext; 
wire [31:0] qa, qb; 
wire [1:0] fwda, fwdb; 
wire [15:0] s16 = {16{sext & inst[15]}};
wire [31:0] dis = {dimm[29:0],2'b00}; 
wire rsrtequ = ~|(a^b); 
pipeidcu cu (mwreg,mrn,ern,ewreg,em2reg,mm2reg,rsrtequ,func,op,rs,rt,wreg,m2reg,wmem,aluc,regrt,aluimm,fwda,fwdb,nostall,sext,pcsrc,shift,jal);
regfile r_f (rs,rt,wdi,wrn,wwreg,~clk,clrn,qa,qb); 
mux2x5 d_r (rd,rt,regrt,rn); 
mux4x32 s_a (qa,ealu,malu,mmo,fwda,a); 
mux4x32 s_b (qb,ealu,malu,mmo,fwdb,b); 
cla32 b_adr (dpc4,dis,1'b0,bpc); 
assign dimm = {s16,imm}; 
assign jpc = {dpc4[31:28],addr,2'b00}; 
endmodule